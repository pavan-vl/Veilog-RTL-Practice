//Designed by Pavan V L
module atm_sys();

endmodule