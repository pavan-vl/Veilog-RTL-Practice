//Designed by Pavan V L
module ele_ctrl();
endmodule