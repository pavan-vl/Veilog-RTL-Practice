//Designed by Pavan V L
module wash_mach();

endmodule