//Designed by Pavan V L
module dig_lock_sys();

endmodule