//Designed by Pavan V L
module euc_gcd(  );
