//Designed by Pavan V L
module rem_sys();

endmodule