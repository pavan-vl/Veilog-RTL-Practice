//Designed by Pavan V L
module feistel_ciph();
endmodule