//Designed by Pavan V L
module tmp_ctrl();
endmodule