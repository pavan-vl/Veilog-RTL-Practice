//Designed by Pavan V L
module ser_int();



endmodule