//Designed by Pavan V L
module irri_sys();

endmodule