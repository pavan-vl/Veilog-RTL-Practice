module uart_tb;
reg clk=0;
reg start=0;
reg [7:0]txin;
wire [7:0]rxout;
wire rxdone,txdone;
     
wire tx2rx;
integer i=0;
       
uart uart_inst(clk,start,tx2rx,txin,tx2rx,rxdone,txdone,rxout);
     
initial begin
start=1;
for(i=0;i<10;i=i+1) begin
txin=$urandom_range(10,200);
@(posedge rxdone);
@(posedge txdone);
end
$finish; 
end
     
always #5 clk = ~clk;
     
endmodule
